`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 18.11.2024 16:13:19
// Design Name: 
// Module Name: MEMORY
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MAIN_MEM (input [15 : 0] addr,din,
output reg [15 : 0] memout,
input rw,
input clk,
input en,
input rst
);

//reg [15 : 0] ram [0 : 1<<13];  //2^13 memory addresses
reg[15 : 0] ram[0 : 1<<8];
//always @(posedge rst) begin   //write your memory here

//end
//always @(posedge rst) begin



always @(*) begin
//if(en) memout <= ram[addr[12 : 0]];
if(en) memout <= ram[addr[7 : 0]]; /// lets use 256 X 16 bits memory
else memout <= 16'b0000_0000_0000_0000;
end
always @(posedge clk or posedge rst) begin
if(rst) begin
ram[0] = 16'b1100_000_000_000_000  ; //mov r0 #0
ram[1] = 16'b0000_0000_0000_0000;
ram[2] = 16'b1100_000_001_000_000  ; //mov r1 #1 
ram[3] = 16'b0000_0000_0000_0001;
ram[4] = 16'b1100_000_011_000_000  ; //mov r3 #10  
ram[5] = 16'b0000_0000_0000_1010;
ram[6] = 16'b1100_000_111_000_000  ; //mov r7 #12
ram[7] = 16'b0000_0000_0000_1100;
ram[8] = 16'b1100_000_100_000_000  ; //mov r4 #2      
ram[9] = 16'b0000_0000_0000_0010;
ram[10] = 16'b1100_000_101_000_000  ; //mov r5 #1   
ram[11] = 16'b0000_0000_0000_0001;
ram[12] = 16'b0001_000_010_001_000  ; //add r2 r1 r0
ram[14] = 16'b1011_000_000_001_000  ; //mov r0 r1
ram[16] = 16'b1011_000_001_010_000  ; //mov r1 r2
ram[18] = 16'b0001_000_100_100_101  ; //add r4 r4 r5    
ram[20] = 16'b1001_000_000_100_011  ; //cmp r4 r3   
ram[22] = 16'b1010_101_000_000_000  ; //skip ge 
ram[24] = 16'b0110_000_111_000_000  ; //jmp r7
ram[26] = 16'b1111_000_000_000_000  ; //halt
end
else if(en)begin
if(rw) ram[addr[7 : 0]] <= din;
end
end
endmodule

module CON_MEM (input [7 : 0] addr,
output reg [15 : 0] memout,
input en,
input rst
);



reg [15 : 0] ram [0 : 1<<8];  //2^13 memory addresses

always @(posedge rst)begin
ram[8'b00000000]=16'b0000000000001000 ;
ram[8'b00000001]=16'b0000100000000100 ;
ram[8'b00010000]=16'b0001000010001000 ;
ram[8'b00010001]=16'b0011100010010000 ;
ram[8'b00010010]=16'b0100000000000000 ;
ram[8'b00100000]=16'b0001100100001000 ;
ram[8'b00100001]=16'b0011100100010000 ;
ram[8'b00100010]=16'b0100000000000000 ;
ram[8'b00110000]=16'b0010100110001000 ;
ram[8'b00110001]=16'b0011100110010000 ;
ram[8'b00110010]=16'b0100000000000000 ;
ram[8'b01000000]=16'b0010001000001000 ;
ram[8'b01000001]=16'b0011101000010000 ;
ram[8'b01000010]=16'b0100000000000000 ;
ram[8'b01010000]=16'b0011001010001000 ;
ram[8'b01010001]=16'b0011101010010000 ;
ram[8'b01010010]=16'b0100000000000000 ;
ram[8'b01100000]=16'b0100101100001000 ;
ram[8'b01100001]=16'b0101001100010000 ;
ram[8'b01100010]=16'b1011000000000000 ;
ram[8'b10100000]=16'b0111000000000000 ;
ram[8'b10010000]=16'b1100000000000000 ;
ram[8'b10110000]=16'b1011110110001000 ;
ram[8'b10110001]=16'b0100000000000000 ;
ram[8'b11000000]=16'b0101111000001000 ;
ram[8'b11000001]=16'b0110111000010000 ;
ram[8'b11000010]=16'b0100000000000000 ;
ram[8'b11010000]=16'b1010011010001000 ;
ram[8'b11010001]=16'b0100000000000000 ;
ram[8'b11100000]=16'b0100111100001000 ;
ram[8'b11100001]=16'b1010100000000000 ;
ram[8'b11110000]=16'b1000011110000000 ;
ram[8'b01110000]=16'b1011101110001000 ;
ram[8'b01110001]=16'b0101001110010000 ;
ram[8'b01110010]=16'b0110101110011000 ;
ram[8'b01110011]=16'b0100000000000000 ;
ram[8'b10000000]=16'b1011110000001000 ;
ram[8'b10000001]=16'b0101010000010000 ;
ram[8'b10000010]=16'b0100110000011000 ;
ram[8'b10000011]=16'b0110000000000000 ;
end

always @(*) begin
if(en) memout <= ram[addr];
end


endmodule





